module NAME3(
  // Write your IO Port Declarations here
  output bit[3:0] y
);  
  assign y = 4'b1111;
  bit a;
  assign a = 1'b0;
endmodule