module not_not_gate(
  input bit a,
  output bit y
  
);  
  // Write your Assignments here
  not_gate n1 (.a(a), .y(y));
  
  
  
endmodule