module NAME(
  input bit a,
  output bit y
  
);  
  // Write your Assignments here
  assign y = ~a; 
  
  
  
endmodule