module not_gate(
  // Write your IO Port Declarations here
  input bit a,
  output bit y
  
);  
  // Write your Assignments here
  assign y = ~a;
  
  
  
endmodule