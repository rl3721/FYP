module NAME2(
  // Write your IO Port Declarations here
  input bit [1:0] a,
  output bit [1:0] y
  
);  
  // Write your Assignments here
  assign y = a;
  
  
  
endmodule